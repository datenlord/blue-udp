
`define SIM_SPEED_UP
