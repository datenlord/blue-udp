import UdpReceiver::*;

(* synthesize *)
module mkTestUdpReceiver();
    UdpReceiver udpReceiver <- mkUdpReceiver;
endmodule