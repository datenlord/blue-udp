`define BSV_POSITIVE_RESET

`define SIM_SPEED_UP