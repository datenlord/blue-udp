
// LRH(64 bits of 1's) + IP Frame
// TTL=1's TOS = 1's Header Checksum = 1's
// UDP Checksum = 1's


// Total Length of IP Frame contains ICRC field
// Total Length of UDP Frame contains ICRC field

// Resv8a field?
// CRC Verification in RX ?











